module hi();
// input and output
endmodule