module hi();

endmodule