module TDC(
	input wire clk,
	input wire pulse1,
	input wire pulse2,
	output reg [7:0] START_END_INTERVAL // [7] START , [6] END, [5:0] INTERVAL 
);

endmodule

