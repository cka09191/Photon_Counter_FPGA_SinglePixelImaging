module TDC(
	input wire clk,
	input wire pulse1,
	input wire pulse2,
	output reg START,
	output reg END,
	output reg [5:0] INTERVAL,
	output reg data_arrived
);

endmodule

