library verilog;
use verilog.vl_types.all;
entity DataMemory is
    port(
        clk             : in     vl_logic;
        RD              : in     vl_logic;
        DMD_sig         : in     vl_logic;
        data_in         : in     vl_logic_vector(15 downto 0);
        rxValid         : in     vl_logic;
        data_out        : out    vl_logic_vector(15 downto 0)
    );
end DataMemory;
