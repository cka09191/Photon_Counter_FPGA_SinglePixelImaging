module Pulse_Shaper(
	input wire clk,
	input wire channel,
	output wire pulse
);

endmodule
