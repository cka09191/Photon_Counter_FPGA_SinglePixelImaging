library verilog;
use verilog.vl_types.all;
entity tb_counter is
end tb_counter;
