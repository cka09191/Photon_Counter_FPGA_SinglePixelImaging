module Command(
	input wire clk,
	input wire [8191:0] rx,
	output reg [1:0] Command
);

endmodule